// Copyright 2021 The CFU-Playground Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.



module Vfu (
  input              cmd_valid,
  output             cmd_ready,
  input     [31:0]   cmd_payload_instruction,
  input     [31:0]   cmd_payload_inputs_0,
  input     [31:0]   cmd_payload_inputs_1,
  input     [2:0]    cmd_payload_rounding,
  output             rsp_valid,
  input              rsp_ready,
  output      [31:0] rsp_payload_output,

  input              reset,
  input              clk
);

  // Trivial handshaking for a combinational CFU
  assign rsp_valid = cmd_valid;
  assign cmd_ready = rsp_ready;

  //
  // select output -- note that we're not fully decoding the 3 function_id bits
  //
  assign rsp_payload_output = cmd_payload_instruction[0] ? 
                                cmd_payload_inputs_1 :
                                cmd_payload_inputs_0 ;


endmodule
